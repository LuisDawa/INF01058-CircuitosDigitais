library verilog;
use verilog.vl_types.all;
entity SCLA_vlg_vec_tst is
end SCLA_vlg_vec_tst;
