library verilog;
use verilog.vl_types.all;
entity lab071_vlg_vec_tst is
end lab071_vlg_vec_tst;
