library verilog;
use verilog.vl_types.all;
entity RCA8bits_vlg_vec_tst is
end RCA8bits_vlg_vec_tst;
