library verilog;
use verilog.vl_types.all;
entity LAB06_vlg_vec_tst is
end LAB06_vlg_vec_tst;
