library verilog;
use verilog.vl_types.all;
entity RCA_vlg_vec_tst is
end RCA_vlg_vec_tst;
