library verilog;
use verilog.vl_types.all;
entity ArithmeticUnit_vlg_vec_tst is
end ArithmeticUnit_vlg_vec_tst;
