library verilog;
use verilog.vl_types.all;
entity lab071 is
    port(
        Q               : out    vl_logic;
        clk             : in     vl_logic
    );
end lab071;
