library verilog;
use verilog.vl_types.all;
entity RCA16bits_vlg_vec_tst is
end RCA16bits_vlg_vec_tst;
