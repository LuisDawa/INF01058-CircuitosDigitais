library verilog;
use verilog.vl_types.all;
entity RCA4bits_vlg_vec_tst is
end RCA4bits_vlg_vec_tst;
