library verilog;
use verilog.vl_types.all;
entity LAB06_vlg_check_tst is
    port(
        A_D             : in     vl_logic;
        B_D             : in     vl_logic;
        C_D             : in     vl_logic;
        D_D             : in     vl_logic;
        E_D             : in     vl_logic;
        F_D             : in     vl_logic;
        G_D             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end LAB06_vlg_check_tst;
