library verilog;
use verilog.vl_types.all;
entity encod_vlg_vec_tst is
end encod_vlg_vec_tst;
