library verilog;
use verilog.vl_types.all;
entity LAB08_vlg_vec_tst is
end LAB08_vlg_vec_tst;
